// system.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module system (
		input  wire        clk_clk,                                            //                              clk.clk
		input  wire [4:0]  pll_0_cntsel_cntsel,                                //                     pll_0_cntsel.cntsel
		output wire        pll_0_outclk0_clk,                                  //                    pll_0_outclk0.clk
		output wire        pll_0_phase_done_phase_done,                        //                 pll_0_phase_done.phase_done
		input  wire        pll_0_phase_en_phase_en,                            //                   pll_0_phase_en.phase_en
		output wire [63:0] pll_0_reconfig_from_pll_reconfig_from_pll,          //          pll_0_reconfig_from_pll.reconfig_from_pll
		input  wire [63:0] pll_0_reconfig_to_pll_reconfig_to_pll,              //            pll_0_reconfig_to_pll.reconfig_to_pll
		input  wire        pll_0_updn_updn,                                    //                       pll_0_updn.updn
		output wire        pll_reconfig_0_mgmt_avalon_slave_waitrequest,       // pll_reconfig_0_mgmt_avalon_slave.waitrequest
		input  wire        pll_reconfig_0_mgmt_avalon_slave_read,              //                                 .read
		input  wire        pll_reconfig_0_mgmt_avalon_slave_write,             //                                 .write
		output wire [31:0] pll_reconfig_0_mgmt_avalon_slave_readdata,          //                                 .readdata
		input  wire [5:0]  pll_reconfig_0_mgmt_avalon_slave_address,           //                                 .address
		input  wire [31:0] pll_reconfig_0_mgmt_avalon_slave_writedata,         //                                 .writedata
		input  wire [63:0] pll_reconfig_0_reconfig_from_pll_reconfig_from_pll, // pll_reconfig_0_reconfig_from_pll.reconfig_from_pll
		output wire [63:0] pll_reconfig_0_reconfig_to_pll_reconfig_to_pll,     //   pll_reconfig_0_reconfig_to_pll.reconfig_to_pll
		input  wire        reset_reset_n                                       //                            reset.reset_n
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> pll_reconfig_0:mgmt_reset

	system_pll_0 pll_0 (
		.refclk            (clk_clk),                                   //            refclk.clk
		.rst               (~reset_reset_n),                            //             reset.reset
		.outclk_0          (pll_0_outclk0_clk),                         //           outclk0.clk
		.phase_en          (pll_0_phase_en_phase_en),                   //          phase_en.phase_en
		.updn              (pll_0_updn_updn),                           //              updn.updn
		.cntsel            (pll_0_cntsel_cntsel),                       //            cntsel.cntsel
		.phase_done        (pll_0_phase_done_phase_done),               //        phase_done.phase_done
		.reconfig_to_pll   (pll_0_reconfig_to_pll_reconfig_to_pll),     //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_0_reconfig_from_pll_reconfig_from_pll), // reconfig_from_pll.reconfig_from_pll
		.locked            ()                                           //       (terminated)
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64)
	) pll_reconfig_0 (
		.mgmt_clk          (clk_clk),                                            //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_reset_out_reset),                     //        mgmt_reset.reset
		.mgmt_waitrequest  (pll_reconfig_0_mgmt_avalon_slave_waitrequest),       // mgmt_avalon_slave.waitrequest
		.mgmt_read         (pll_reconfig_0_mgmt_avalon_slave_read),              //                  .read
		.mgmt_write        (pll_reconfig_0_mgmt_avalon_slave_write),             //                  .write
		.mgmt_readdata     (pll_reconfig_0_mgmt_avalon_slave_readdata),          //                  .readdata
		.mgmt_address      (pll_reconfig_0_mgmt_avalon_slave_address),           //                  .address
		.mgmt_writedata    (pll_reconfig_0_mgmt_avalon_slave_writedata),         //                  .writedata
		.reconfig_to_pll   (pll_reconfig_0_reconfig_to_pll_reconfig_to_pll),     //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_reconfig_0_reconfig_from_pll_reconfig_from_pll), // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                             //       (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
